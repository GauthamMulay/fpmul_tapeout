magic
tech sky130A
magscale 1 2
timestamp 1700845427
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 934 2128 558808 349840
<< metal2 >>
rect 279974 0 280030 800
<< obsm2 >>
rect 938 856 558422 349829
rect 938 800 279918 856
rect 280086 800 558422 856
<< metal3 >>
rect 0 342184 800 342304
rect 559200 338920 560000 339040
rect 0 323688 800 323808
rect 559200 317160 560000 317280
rect 0 305192 800 305312
rect 559200 295400 560000 295520
rect 0 286696 800 286816
rect 559200 273640 560000 273760
rect 0 268200 800 268320
rect 559200 251880 560000 252000
rect 0 249704 800 249824
rect 0 231208 800 231328
rect 559200 230120 560000 230240
rect 0 212712 800 212832
rect 559200 208360 560000 208480
rect 0 194216 800 194336
rect 559200 186600 560000 186720
rect 0 175720 800 175840
rect 559200 164840 560000 164960
rect 0 157224 800 157344
rect 559200 143080 560000 143200
rect 0 138728 800 138848
rect 559200 121320 560000 121440
rect 0 120232 800 120352
rect 0 101736 800 101856
rect 559200 99560 560000 99680
rect 0 83240 800 83360
rect 559200 77800 560000 77920
rect 0 64744 800 64864
rect 559200 56040 560000 56160
rect 0 46248 800 46368
rect 559200 34280 560000 34400
rect 0 27752 800 27872
rect 559200 12520 560000 12640
rect 0 9256 800 9376
<< obsm3 >>
rect 800 342384 559200 349825
rect 880 342104 559200 342384
rect 800 339120 559200 342104
rect 800 338840 559120 339120
rect 800 323888 559200 338840
rect 880 323608 559200 323888
rect 800 317360 559200 323608
rect 800 317080 559120 317360
rect 800 305392 559200 317080
rect 880 305112 559200 305392
rect 800 295600 559200 305112
rect 800 295320 559120 295600
rect 800 286896 559200 295320
rect 880 286616 559200 286896
rect 800 273840 559200 286616
rect 800 273560 559120 273840
rect 800 268400 559200 273560
rect 880 268120 559200 268400
rect 800 252080 559200 268120
rect 800 251800 559120 252080
rect 800 249904 559200 251800
rect 880 249624 559200 249904
rect 800 231408 559200 249624
rect 880 231128 559200 231408
rect 800 230320 559200 231128
rect 800 230040 559120 230320
rect 800 212912 559200 230040
rect 880 212632 559200 212912
rect 800 208560 559200 212632
rect 800 208280 559120 208560
rect 800 194416 559200 208280
rect 880 194136 559200 194416
rect 800 186800 559200 194136
rect 800 186520 559120 186800
rect 800 175920 559200 186520
rect 880 175640 559200 175920
rect 800 165040 559200 175640
rect 800 164760 559120 165040
rect 800 157424 559200 164760
rect 880 157144 559200 157424
rect 800 143280 559200 157144
rect 800 143000 559120 143280
rect 800 138928 559200 143000
rect 880 138648 559200 138928
rect 800 121520 559200 138648
rect 800 121240 559120 121520
rect 800 120432 559200 121240
rect 880 120152 559200 120432
rect 800 101936 559200 120152
rect 880 101656 559200 101936
rect 800 99760 559200 101656
rect 800 99480 559120 99760
rect 800 83440 559200 99480
rect 880 83160 559200 83440
rect 800 78000 559200 83160
rect 800 77720 559120 78000
rect 800 64944 559200 77720
rect 880 64664 559200 64944
rect 800 56240 559200 64664
rect 800 55960 559120 56240
rect 800 46448 559200 55960
rect 880 46168 559200 46448
rect 800 34480 559200 46168
rect 800 34200 559120 34480
rect 800 27952 559200 34200
rect 880 27672 559200 27952
rect 800 12720 559200 27672
rect 800 12440 559120 12720
rect 800 9456 559200 12440
rect 880 9176 559200 9456
rect 800 2143 559200 9176
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< labels >>
rlabel metal3 s 559200 12520 560000 12640 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 268200 800 268320 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 231208 800 231328 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 194216 800 194336 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 175720 800 175840 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 157224 800 157344 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 138728 800 138848 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 120232 800 120352 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 0 101736 800 101856 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 559200 56040 560000 56160 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 559200 99560 560000 99680 6 io_in[2]
port 16 nsew signal input
rlabel metal3 s 559200 143080 560000 143200 6 io_in[3]
port 17 nsew signal input
rlabel metal3 s 559200 186600 560000 186720 6 io_in[4]
port 18 nsew signal input
rlabel metal3 s 559200 230120 560000 230240 6 io_in[5]
port 19 nsew signal input
rlabel metal3 s 559200 273640 560000 273760 6 io_in[6]
port 20 nsew signal input
rlabel metal3 s 559200 317160 560000 317280 6 io_in[7]
port 21 nsew signal input
rlabel metal3 s 0 342184 800 342304 6 io_in[8]
port 22 nsew signal input
rlabel metal3 s 0 305192 800 305312 6 io_in[9]
port 23 nsew signal input
rlabel metal3 s 559200 34280 560000 34400 6 io_out[0]
port 24 nsew signal output
rlabel metal3 s 0 249704 800 249824 6 io_out[10]
port 25 nsew signal output
rlabel metal3 s 0 212712 800 212832 6 io_out[11]
port 26 nsew signal output
rlabel metal3 s 559200 77800 560000 77920 6 io_out[1]
port 27 nsew signal output
rlabel metal3 s 559200 121320 560000 121440 6 io_out[2]
port 28 nsew signal output
rlabel metal3 s 559200 164840 560000 164960 6 io_out[3]
port 29 nsew signal output
rlabel metal3 s 559200 208360 560000 208480 6 io_out[4]
port 30 nsew signal output
rlabel metal3 s 559200 251880 560000 252000 6 io_out[5]
port 31 nsew signal output
rlabel metal3 s 559200 295400 560000 295520 6 io_out[6]
port 32 nsew signal output
rlabel metal3 s 559200 338920 560000 339040 6 io_out[7]
port 33 nsew signal output
rlabel metal3 s 0 323688 800 323808 6 io_out[8]
port 34 nsew signal output
rlabel metal3 s 0 286696 800 286816 6 io_out[9]
port 35 nsew signal output
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 37 nsew ground bidirectional
rlabel metal2 s 279974 0 280030 800 6 wb_clk_i
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 52765054
string GDS_FILE /home/kiran/special_topic_asics/fpmul_tapeout/openlane/user_proj_example/runs/23_11_24_22_18/results/signoff/user_proj_example.magic.gds
string GDS_START 433266
<< end >>

